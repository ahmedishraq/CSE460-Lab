module inverter_lab06(A,Y);

	input A;
	output Y;

	not(Y,A);

endmodule